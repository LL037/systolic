// mac_array.v
// MAC array module
// Composes multiple MAC units into an array
// Inputs:
//  - clk: clock signal
//  - rst: reset signal
//  - valid_ctrl: control signals for each MAC unit
//  - clear: clear signals for each MAC unit
// - valid_weight_in: weight valid signals for each MAC unit
//  - a_in: single activation input (flows through the array)
//  - w_0, w_1, w_2, w_3: weight inputs for each MAC unit
// Outputs:
// - acc_out_0, acc_out_1, acc_out_2, acc_out_3: accumulator outputs from each MAC unit
//  - valid_out: valid output signals from each MAC unit


module mac_array #(
    parameter W      = 8,  
    parameter ACC_W  = 16,
    parameter N_MACS = 4
)(
    input  wire                    clk,
    input  wire                    rst,

    input  wire [3*N_MACS-1:0]     valid_ctrl,
 
    input  wire [N_MACS-1:0]       clear, 
    input  wire [N_MACS-1:0]       valid_weight_in,
     
    // Single activation input (flows through the array)
    input  wire signed [ACC_W-1:0]     a_in,
    
    // Weight inputs for each MAC
    input  wire signed [ACC_W-1:0]     w_0,        // Weight for MAC 0
    input  wire signed [ACC_W-1:0]     w_1,        // Weight for MAC 1
    input  wire signed [ACC_W-1:0]     w_2,        // Weight for MAC 2
    input  wire signed [ACC_W-1:0]     w_3,        // Weight for MAC 3
    
    // Final outputs
    output wire signed [ACC_W-1:0] acc_out_0,
    output wire signed [ACC_W-1:0] acc_out_1,
    output wire signed [ACC_W-1:0] acc_out_2,
    output wire signed [ACC_W-1:0] acc_out_3,
    output wire [N_MACS-1:0]       valid_out
);

    wire signed [ACC_W-1:0]     a_out_0_1;
    wire signed [ACC_W-1:0]     a_out_0_1_1;

    wire signed [ACC_W-1:0]     a_out_1_0;  
    wire signed [ACC_W-1:0]     a_out_2_3;  
    wire signed [ACC_W-1:0]     a_out_3_2; 
    wire [2:0] valid_ctrl_0;
    wire [2:0] valid_ctrl_1;
    wire [2:0] valid_ctrl_2;
    wire [2:0] valid_ctrl_3;



    assign valid_ctrl_0 = valid_ctrl[2:0];
    assign valid_ctrl_1 = valid_ctrl[5:3];
    assign valid_ctrl_2 = valid_ctrl[8:6];
    assign valid_ctrl_3 = valid_ctrl[11:9];


    // MAC 0 (top-left)
    mac #(
        .W(W),
        .ACC_W(ACC_W)
    ) mac_0 (
        .clk(clk),
        .rst(rst),
        .acc_sel(3'b000),
        .valid_ctrl(valid_ctrl_0),
        .weight_valid_in(valid_weight_in[0]),
        .clear(clear[0]),
        .a_in_0(a_in),
        .a_in_1(acc_out_2),
        .a_in_2(a_out_1_0),              
        .weight(w_0),               
        .acc_out(acc_out_0),
        .valid_out(valid_out[0]),
        .a_out_0(a_out_0_1),
        .a_out_1(a_out_0_1_1),
        .a_out_2()        
    );

    // MAC 1 (top-right)
    mac #(
        .W(W),
        .ACC_W(ACC_W)
    ) mac_1 (
        .clk(clk),
        .rst(rst),
        .acc_sel(3'b000),
        .valid_ctrl(valid_ctrl_1),
        .weight_valid_in(valid_weight_in[1]),
        .clear(clear[1]),
        .a_in_0(a_out_0_1),
        .a_in_1(a_out_0_1_1),   
        .a_in_2(acc_out_3),            
        .weight(w_1),               
        .acc_out(acc_out_1),
        .valid_out(valid_out[1]),
        .a_out_0(),
        .a_out_1(),
        .a_out_2(a_out_1_0)        
    );

    // MAC 2 (bottom-left)
    mac #(
        .W(W),
        .ACC_W(ACC_W)
    ) mac_2 (
        .clk(clk),
        .rst(rst),
        .acc_sel(3'b000),
        .valid_ctrl(valid_ctrl_2),
        .weight_valid_in(valid_weight_in[2]),
        .clear(clear[2]),
        .a_in_0(acc_out_0),
        .a_in_1(a_out_3_2),
        .a_in_2(),                
        .weight(w_2),               
        .acc_out(acc_out_2),
        .valid_out(valid_out[2]),
        .a_out_0(a_out_2_3),
        .a_out_1(), 
        .a_out_2()        
       
    );
    // MAC 3 (bottom-right)
    mac #(
        .W(W),
        .ACC_W(ACC_W)
    ) mac_3 (
        .clk(clk),
        .rst(rst),
        .acc_sel(3'b000),
        .valid_ctrl(valid_ctrl_3),
        .weight_valid_in(valid_weight_in[3]),
        .clear(clear[3]),
        .a_in_0(acc_out_1),
        .a_in_1(a_out_2_3), 
        .a_in_2(),             
        .weight(w_3),               
        .acc_out(acc_out_3),
        .valid_out(valid_out[3]),
        .a_out_0(a_out_3_2),
        .a_out_1(),  
        .a_out_2()        

    );

endmodule
